LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY top_level_timer IS
    PORT (
        CLOCK_50 : IN STD_LOGIC;
        SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
        KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
        LEDR : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
        HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
        HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE Behavioral OF top_level_timer IS

    -- === Clock division ===
    SIGNAL clk_divider : unsigned(25 DOWNTO 0) := (OTHERS => '0');
    SIGNAL one_hz_clk : STD_LOGIC := '0';
    SIGNAL tick_1hz : STD_LOGIC := '0';

    -- === Timer I/O Signals ===
    SIGNAL Q_sec_ones : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL Q_sec_tens : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL Q_min_ones : STD_LOGIC_VECTOR(3 DOWNTO 0);

    -- === Control ===
    SIGNAL Enable : STD_LOGIC := '0';
    SIGNAL Reset : STD_LOGIC := '0';
    SIGNAL initial_switch_value : STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');

    SIGNAL send_to_reset_1 : STD_LOGIC := '0';

    SIGNAL send_to_Enable_1 : STD_LOGIC := '0';
    SIGNAL send_to_Enable_2 : STD_LOGIC := '1';


    -- Captured values (capped)
    signal target_sec_ones  : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
    signal target_sec_tens  : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
    signal target_min_ones  : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

    -- === Component declarations ===
    COMPONENT three_digit_timer
        PORT (
            Clk : IN STD_LOGIC;
            Reset : IN STD_LOGIC;
            Enable : IN STD_LOGIC;
            Min_ones : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            Sec_tens : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            Sec_ones : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT BCD_to_SevenSeg
        PORT (
            BCD_digit : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            SevenSeg_out : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
        );
    END COMPONENT;

BEGIN

    -- === Button press logic ===
    PROCESS (CLOCK_50)
    variable sw_ones  : unsigned(3 downto 0);
    variable sw_tens  : unsigned(3 downto 0);
    variable sw_mins  : unsigned(1 downto 0);
BEGIN
    IF rising_edge(CLOCK_50) THEN
        IF KEY(0) = '0' THEN  -- Button pressed (active-low)

            -- Store full raw switch value
            initial_switch_value <= SW;

            -- === CAP AND STORE EACH SECTION ===
            sw_ones := unsigned(SW(3 downto 0));
            IF sw_ones > 9 THEN
                target_sec_ones <= "1001";  -- 9
            ELSE
                target_sec_ones <= std_logic_vector(sw_ones);
            END IF;

            sw_tens := unsigned(SW(7 downto 4));
            IF sw_tens > 5 THEN
                target_sec_tens <= "0101";  -- 5
            ELSE
                target_sec_tens <= std_logic_vector(sw_tens);
            END IF;

            sw_mins := unsigned(SW(9 downto 8));
            IF sw_mins > 3 THEN
                target_min_ones <= "0011";  -- 3
            ELSE
                target_min_ones <= "00" & std_logic_vector(sw_mins);  -- Now it's 4 bits
            END IF;

            -- Trigger timer reset & enable
            send_to_Enable_1 <= '1';
            send_to_reset_1 <= '1';

        ELSE
            send_to_reset_1 <= '0';
        END IF;
    END IF;
END PROCESS;
    -- === Clock Divider ===
    PROCESS (CLOCK_50)
    BEGIN
        IF rising_edge(CLOCK_50) THEN
            IF clk_divider = 4_999_999 THEN -- 50 MHz ÷ 50M = 1Hz (original is 49_999_999)
                clk_divider <= (OTHERS => '0');
                one_hz_clk <= NOT one_hz_clk;
                tick_1hz <= '1';
            ELSE
                clk_divider <= clk_divider + 1;
                tick_1hz <= '0';
            END IF;
        END IF;
    END PROCESS;

    -- === Timer Instance ===
    timer_inst : three_digit_timer
    PORT MAP(
        Clk => tick_1hz,
        Reset => Reset,
        Enable => Enable,
        Min_ones => Q_min_ones,
        Sec_tens => Q_sec_tens,
        Sec_ones => Q_sec_ones
    );

    -- === Seven Segment Display ===
    seg0 : BCD_to_SevenSeg
    PORT MAP(
        BCD_digit => Q_sec_ones,
        SevenSeg_out => HEX0
    );

    seg1 : BCD_to_SevenSeg
    PORT MAP(
        BCD_digit => Q_sec_tens,
        SevenSeg_out => HEX1
    );

    seg2 : BCD_to_SevenSeg
    PORT MAP(
        BCD_digit => Q_min_ones,
        SevenSeg_out => HEX2
    );



    -- Stop counting when the timer reaches the stored value
    PROCESS (CLOCK_50)
    BEGIN
        IF rising_edge(CLOCK_50) THEN
            IF Enable = '1' THEN
                IF Q_min_ones = target_min_ones AND
                Q_sec_tens = target_sec_tens AND
                Q_sec_ones = target_sec_ones THEN
                    send_to_Enable_2 <= '0';  -- Stop counting
                END IF;
            ELSE
                send_to_Enable_2 <= '1';  -- Resume counting
            END IF;
        END IF;
    END PROCESS;

    Reset <= send_to_reset_1;
    Enable <= send_to_Enable_1 and send_to_Enable_2;

    -- === Debug LED ===
    LEDR(0) <= Enable;
    LEDR(1) <= Reset;

END ARCHITECTURE;